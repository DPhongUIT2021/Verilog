library verilog;
use verilog.vl_types.all;
entity Register8bitBasic_vlg_vec_tst is
end Register8bitBasic_vlg_vec_tst;
