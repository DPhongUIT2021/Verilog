library verilog;
use verilog.vl_types.all;
entity Adder8Bit_vlg_vec_tst is
end Adder8Bit_vlg_vec_tst;
