library verilog;
use verilog.vl_types.all;
entity ControlFunctionSharing_vlg_vec_tst is
end ControlFunctionSharing_vlg_vec_tst;
