library verilog;
use verilog.vl_types.all;
entity Decode_vlg_vec_tst is
end Decode_vlg_vec_tst;
