library verilog;
use verilog.vl_types.all;
entity Max_vlg_vec_tst is
end Max_vlg_vec_tst;
