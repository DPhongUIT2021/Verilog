library verilog;
use verilog.vl_types.all;
entity Decode4To10_vlg_vec_tst is
end Decode4To10_vlg_vec_tst;
