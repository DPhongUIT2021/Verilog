library verilog;
use verilog.vl_types.all;
entity RegisterSharingDatapath_vlg_vec_tst is
end RegisterSharingDatapath_vlg_vec_tst;
