library verilog;
use verilog.vl_types.all;
entity Adder16Bit_vlg_vec_tst is
end Adder16Bit_vlg_vec_tst;
