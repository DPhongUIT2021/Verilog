library verilog;
use verilog.vl_types.all;
entity OneRegister16bit_vlg_vec_tst is
end OneRegister16bit_vlg_vec_tst;
