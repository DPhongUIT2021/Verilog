library verilog;
use verilog.vl_types.all;
entity AbsMax_vlg_vec_tst is
end AbsMax_vlg_vec_tst;
