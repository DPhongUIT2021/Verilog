library verilog;
use verilog.vl_types.all;
entity ShiftRight3bit_vlg_vec_tst is
end ShiftRight3bit_vlg_vec_tst;
