library verilog;
use verilog.vl_types.all;
entity ShiftRight1bit_vlg_vec_tst is
end ShiftRight1bit_vlg_vec_tst;
