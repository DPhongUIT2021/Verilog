library verilog;
use verilog.vl_types.all;
entity Mux4To1Shift_vlg_check_tst is
    port(
        O               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Mux4To1Shift_vlg_check_tst;
