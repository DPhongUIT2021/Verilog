library verilog;
use verilog.vl_types.all;
entity AddSub16bit_vlg_vec_tst is
end AddSub16bit_vlg_vec_tst;
