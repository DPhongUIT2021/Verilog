library verilog;
use verilog.vl_types.all;
entity MinAbsAddSub_vlg_vec_tst is
end MinAbsAddSub_vlg_vec_tst;
