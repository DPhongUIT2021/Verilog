library verilog;
use verilog.vl_types.all;
entity RFC_vlg_vec_tst is
end RFC_vlg_vec_tst;
