
module SRA_Controler_Beha(ctrl_word, In1, In2, reset, clk);
			parameter msb = 15;
			input[msb:0] In1, In2;
			input reset, clk;
			output ctrl_word;
			
endmodule
