library verilog;
use verilog.vl_types.all;
entity Mux4To1Shift_vlg_vec_tst is
end Mux4To1Shift_vlg_vec_tst;
