library verilog;
use verilog.vl_types.all;
entity ShiftRight1_16bit_vlg_vec_tst is
end ShiftRight1_16bit_vlg_vec_tst;
