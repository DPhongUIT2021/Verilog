library verilog;
use verilog.vl_types.all;
entity ShiftRight3_16it_vlg_vec_tst is
end ShiftRight3_16it_vlg_vec_tst;
