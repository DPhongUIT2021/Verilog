library verilog;
use verilog.vl_types.all;
entity Latch16bit_vlg_vec_tst is
end Latch16bit_vlg_vec_tst;
