library verilog;
use verilog.vl_types.all;
entity Mux16Bit_vlg_vec_tst is
end Mux16Bit_vlg_vec_tst;
