library verilog;
use verilog.vl_types.all;
entity AddSubUpdate_vlg_vec_tst is
end AddSubUpdate_vlg_vec_tst;
