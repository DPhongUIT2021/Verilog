library verilog;
use verilog.vl_types.all;
entity Min_vlg_vec_tst is
end Min_vlg_vec_tst;
