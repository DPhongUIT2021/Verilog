library verilog;
use verilog.vl_types.all;
entity FourReg16bit_vlg_vec_tst is
end FourReg16bit_vlg_vec_tst;
