library verilog;
use verilog.vl_types.all;
entity Multi2_vlg_vec_tst is
end Multi2_vlg_vec_tst;
