library verilog;
use verilog.vl_types.all;
entity FourReg16bitTwoInput_vlg_vec_tst is
end FourReg16bitTwoInput_vlg_vec_tst;
