library verilog;
use verilog.vl_types.all;
entity ControlRegisterSharing_vlg_vec_tst is
end ControlRegisterSharing_vlg_vec_tst;
