library verilog;
use verilog.vl_types.all;
entity Mux_4_vlg_vec_tst is
end Mux_4_vlg_vec_tst;
