library verilog;
use verilog.vl_types.all;
entity FunctionUnitSharing_vlg_vec_tst is
end FunctionUnitSharing_vlg_vec_tst;
