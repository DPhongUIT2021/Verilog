library verilog;
use verilog.vl_types.all;
entity Decode2To4_vlg_vec_tst is
end Decode2To4_vlg_vec_tst;
