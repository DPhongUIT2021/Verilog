library verilog;
use verilog.vl_types.all;
entity Multi4_vlg_vec_tst is
end Multi4_vlg_vec_tst;
