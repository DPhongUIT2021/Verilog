library verilog;
use verilog.vl_types.all;
entity Reg16Sharing_vlg_vec_tst is
end Reg16Sharing_vlg_vec_tst;
