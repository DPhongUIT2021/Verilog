

`timescale 1ps/1ps
module tb_SRA_beha();
			

endmodule
