library verilog;
use verilog.vl_types.all;
entity ALULap04_vlg_vec_tst is
end ALULap04_vlg_vec_tst;
