library verilog;
use verilog.vl_types.all;
entity Multi16bit_vlg_vec_tst is
end Multi16bit_vlg_vec_tst;
