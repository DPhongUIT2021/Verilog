library verilog;
use verilog.vl_types.all;
entity RegisterSharing_vlg_vec_tst is
end RegisterSharing_vlg_vec_tst;
