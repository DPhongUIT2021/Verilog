library verilog;
use verilog.vl_types.all;
entity ShiftLeft16bit_vlg_vec_tst is
end ShiftLeft16bit_vlg_vec_tst;
