library verilog;
use verilog.vl_types.all;
entity Latch8bit_vlg_vec_tst is
end Latch8bit_vlg_vec_tst;
