library verilog;
use verilog.vl_types.all;
entity ControlBusSharing_vlg_vec_tst is
end ControlBusSharing_vlg_vec_tst;
