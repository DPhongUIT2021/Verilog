library verilog;
use verilog.vl_types.all;
entity BusSharing_vlg_vec_tst is
end BusSharing_vlg_vec_tst;
