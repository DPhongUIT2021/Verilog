library verilog;
use verilog.vl_types.all;
entity Test1Regiter_vlg_vec_tst is
end Test1Regiter_vlg_vec_tst;
