library verilog;
use verilog.vl_types.all;
entity Mux8Bit_vlg_vec_tst is
end Mux8Bit_vlg_vec_tst;
