library verilog;
use verilog.vl_types.all;
entity Abs_vlg_vec_tst is
end Abs_vlg_vec_tst;
