library verilog;
use verilog.vl_types.all;
entity SRwPL_8bit_vlg_vec_tst is
end SRwPL_8bit_vlg_vec_tst;
