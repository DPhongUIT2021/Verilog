library verilog;
use verilog.vl_types.all;
entity Mux16Bit4To1_vlg_vec_tst is
end Mux16Bit4To1_vlg_vec_tst;
